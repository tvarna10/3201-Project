module round2(clock, round2num1, round2num2, round2num3, round2points, resetswitch, spin, stopkey, fast, slow, testcase);

	input clock;
	input resetswitch;
	input spin;
	input stopkey;
	input fast;
	input slow;
	input testcase;

	// output the generated and selected numbers as well as the points awarded for the round
	// will be used for point addition and number displays
	output reg [7:0] round2points;
	output reg [7:0] round2num1;
	output reg [7:0] round2num2;
	output reg [7:0] round2num3;
	
	// use the numbers generated by the LFSR
	wire [3:0] number1;
	wire [3:0] number2;
	wire [3:0] number3;
	
	// keep track of KEY[1] clicks- keep track each time a number is selected
	wire [3:0] sum;
	reg [3:0] keepspin;
	
	// used for the game speed
	reg speed;

	// instantiate the clocks to determine game speed
   fastspin f1(clock, fastspeed);
	mediumspin m1(clock, moderatespeed);
	slowspin s1(clock, slowspeed);

	// instantiate the LFSR three times to determine the three numbers
	LFSR lfsr1 (speed, resetswitch, number1);
	LFSR lfsr2 (speed, resetswitch, number2);
	LFSR lfsr3 (speed, resetswitch, number3);
	
	fourbitadder f0(keepspin, 4'b0001, 0, sum, carryout);
	
//================================================================================================================//

initial begin
	keepspin <= 4'b0000; // initalize keepspin to 1
end

always @(negedge stopkey) begin // triggered when KEY1 is pressed
	if (!resetswitch) begin // if the reset switch is off
		keepspin <= sum; // keepspin equals sum
	end
	else if (resetswitch) // if reset switch is on
	begin
		keepspin <= 4'b0000; // set keepspin back to 0 -> will allow user to restart the game
	end
end

always @* begin
	case ({fast, slow}) // choose how fast the numbers will spin
		2'b10: speed <= fastspeed; // set speed to fast if switch 2 is up
		2'b01: speed <= slowspeed; // set speed to low if switch 1 is up
		default: speed <= moderatespeed; // set speed to moderate if switch 1 and 2 are down
	endcase
end

always @(posedge speed) begin	

	if (spin) begin

		if (testcase) begin // test cases used to check if point counting and adding worked
								  // can be commented out if not needed
								  // can be removed completely as long as you remove the input from the module and its instances

			round2num1 = 8'b11111000; // set to number 7
			round2num2 = 8'b11111000; // set to number 7
			round2num3 = 8'b11111000; // set to number 7
		
		end
		else begin // if not testcase
		
			if (keepspin == 4'b0011) begin // spin number 1
				
				round2num2 = 8'b11000000; // number 2 initally 0
				round2num3 = 8'b11000000; // number 3 initially 0
			
				case(number1) // will determine the 8 bit value of number 1 based on the random number generated using the LFSR
								  // needs to be 8 bits in order to be used for the display
					4'b1001 : round2num1 = 8'b10010000; // set to number 9
					4'b1000 : round2num1 = 8'b10000000; // set to number 8
					4'b0111 : round2num1 = 8'b11111000; // set to number 7
					4'b0110 : round2num1 = 8'b10000010; // set to number 6
					4'b0101 : round2num1 = 8'b10010010; // set to number 5
					4'b0100 : round2num1 = 8'b10011001; // set to number 4
					4'b0011 : round2num1 = 8'b10110000; // set to number 3
					4'b0010 : round2num1 = 8'b10100100; // set to number 2
					4'b0001 : round2num1 = 8'b11111001; // set to number 1
					4'b0000 : round2num1 = 8'b11000000; // set to number 0
					default : round2num1 = 8'b11000000;
				endcase
			end
			
			if (keepspin == 4'b0100) begin		
				case(number2) // will determine the 8 bit value of number 2 based on the random number generated using the LFSR
								  // needs to be 8 bits in order to be used for the display
					4'b1001 : round2num2= 8'b10010000; // set to number 9
					4'b1000 : round2num2 = 8'b10000000; // set to number 8
					4'b0111 : round2num2 = 8'b11111000; // set to number 7
					4'b0110 : round2num2 = 8'b10000010; // set to number 6
					4'b0101 : round2num2 = 8'b10010010; // set to number 5
					4'b0100 : round2num2 = 8'b10011001; // set to number 4
					4'b0011 : round2num2 = 8'b10110000; // set to number 3
					4'b0010 : round2num2 = 8'b10100100; // set to number 2
					4'b0001 : round2num2 = 8'b11111001; // set to number 1
					4'b0000 : round2num2 = 8'b11000000; // set to number 0
					default : round2num2 = 8'b11000000;
				endcase
			end
			
			if (keepspin == 4'b0101) begin
				case(number3) // will determine the 8 bit value of number 3 based on the random number generated using the LFSR
								  // needs to be 8 bits in order to be used for the display
					4'b1001 : round2num3 = 8'b10010000; // set to number 9
					4'b1000 : round2num3 = 8'b10000000; // set to number 8
					4'b0111 : round2num3 = 8'b11111000; // set to number 7
					4'b0110 : round2num3 = 8'b10000010; // set to number 6
					4'b0101 : round2num3 = 8'b10010010; // set to number 5
					4'b0100 : round2num3 = 8'b10011001; // set to number 4
					4'b0011 : round2num3 = 8'b10110000; // set to number 3
					4'b0010 : round2num3 = 8'b10100100; // set to number 2
					4'b0001 : round2num3 = 8'b11111001; // set to number 1
					4'b0000 : round2num3 = 8'b11000000; // set to number 0
					default : round2num3 = 8'b11000000;
				endcase
			end
		end
	end
end
//================================================================================================================//

always @(posedge speed) begin

	if (resetswitch) begin // if reset switch is on
		round2points <= 8'b00000000; // points automatically go to zero
	end

	else begin // if reset switch is off 
		if (keepspin > 4'b0101) begin // if KEY[1] has been pressed three times (3 numbers have been selected)
					
			// compare the three selected numbers
			if (round2num1 == round2num2 && round2num1 == round2num3) begin // if all the numbers are the same
			
				case(round2num1) // provide a score based off whatever the matched numbers are
					8'b10010000 : round2points = 8'b00011001; // 999 = 25 points
					8'b10000000 : round2points = 8'b00100011; // 888 = 35 points
					8'b11111000 : round2points = 8'b00110010; // 777 = 50 points
					8'b10000010 : round2points = 8'b00100011; // 666 = 35 points
					8'b10010010 : round2points = 8'b00011001; // 555 = 25 points
					8'b10011001 : round2points = 8'b00010100; // 444 = 20 points
					8'b10110000 : round2points = 8'b00001111; // 333 = 15 points
					8'b10100100 : round2points = 8'b00001010; // 222 = 10 points
					8'b11111001 : round2points = 8'b00000101; // 111 = 5 points
					8'b11000000 : round2points = 8'b00000000; // 000 = 0 points
					default : round2points = 8'b00000000;
				endcase
			end
			else begin // if the numbers dont match
				round2points = 8'b00000000; // 0 points are awarded
			end
		end
	end
end

endmodule
